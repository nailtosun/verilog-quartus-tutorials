library verilog;
use verilog.vl_types.all;
entity Mean_vlg_vec_tst is
end Mean_vlg_vec_tst;
