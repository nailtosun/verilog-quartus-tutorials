library verilog;
use verilog.vl_types.all;
entity serial_to_parallel_vlg_vec_tst is
end serial_to_parallel_vlg_vec_tst;
