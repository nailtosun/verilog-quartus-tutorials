library verilog;
use verilog.vl_types.all;
entity frequencyfinder_vlg_vec_tst is
end frequencyfinder_vlg_vec_tst;
